library ieee;
use ieee.std_logic_1164.all;

entity reg_nb is
	
	generic (N: positive := 8);
	port (
		--control inputs
		clk, rst, load: in std_logic;
		--data inputs
		d: in std_logic_vector(N-1 downto 0);
		--data outputs		
		q: out std_logic_vector(N-1 downto 0)
		);
		
end entity;

architecture bhv of reg_nb is

	subtype InternalState is std_logic_vector(N-1 downto 0);
	signal nextState, currentState: InternalState;
	
begin

	-- next-state logic (combinational)
	nextState <= d when load='1' else currentState;
	
	-- memory element (sequential)
	process (clk, rst) is
	begin
		if rst = '1' then
			currentState <= (others => '0'); -- reset state
		elsif rising_edge(clk) then
			currentState <= nextState;
		end if;
	end process;
	
	-- output logic
	q <= currentState;


end bhv;